module mult_1x1 (
    input signed [15:0] a,
    input signed [15:0] b,
    output signed [31:0] out
);

    assign out = a * b;

endmodule
